library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_1164.ALL;

entity clockadjust is
end clockadjust;

architecture Behavioral of clockadjust is

begin


end Behavioral;

